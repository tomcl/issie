module NAME();
bit i, j;

always_comb begin
    i=j;
end

assign j=i;


endmodule