module NAME();
bit i, j;


assign i=j;
assign j=i;


endmodule