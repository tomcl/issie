module NAME();
bit i, j;

always_comb begin
    i=j;
    j=i;
end


endmodule